// -----------------------------------------------------------------------------
// Copyright (c) 1996-2024 All rights reserved
// -----------------------------------------------------------------------------
// Author : wenky
// File : sd_top
// email: wenkyjong1996@gmail.com
// Create : 2024-08-19
// Revise : 
// Functions : 
// 
// -----------------------------------------------------------------------------

module sd_top (
    input   sclk,
    input   rst_n,
    output  sd_clk,
    output 
);
    
endmodule